// qSDRAM_100MHz.v

// Generated using ACDS version 13.1 162 at 2014.04.07.09:24:06

`timescale 1 ps / 1 ps
module qSDRAM_100MHz (
		input  wire        clk_clk,         //   clk.clk
		input  wire        reset_reset_n,   // reset.reset_n
		input  wire [24:0] m_address,       //     m.address
		input  wire [1:0]  m_byteenable_n,  //      .byteenable_n
		input  wire        m_chipselect,    //      .chipselect
		input  wire [15:0] m_writedata,     //      .writedata
		input  wire        m_read_n,        //      .read_n
		input  wire        m_write_n,       //      .write_n
		output wire [15:0] m_readdata,      //      .readdata
		output wire        m_readdatavalid, //      .readdatavalid
		output wire        m_waitrequest,   //      .waitrequest
		output wire [12:0] ram_addr,        //   ram.addr
		output wire [1:0]  ram_ba,          //      .ba
		output wire        ram_cas_n,       //      .cas_n
		output wire        ram_cke,         //      .cke
		output wire        ram_cs_n,        //      .cs_n
		inout  wire [15:0] ram_dq,          //      .dq
		output wire [1:0]  ram_dqm,         //      .dqm
		output wire        ram_ras_n,       //      .ras_n
		output wire        ram_we_n         //      .we_n
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> new_sdram_controller_0:reset_n

	qSDRAM_100MHz_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (clk_clk),                         //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset), // reset.reset_n
		.az_addr        (m_address),                       //    s1.address
		.az_be_n        (m_byteenable_n),                  //      .byteenable_n
		.az_cs          (m_chipselect),                    //      .chipselect
		.az_data        (m_writedata),                     //      .writedata
		.az_rd_n        (m_read_n),                        //      .read_n
		.az_wr_n        (m_write_n),                       //      .write_n
		.za_data        (m_readdata),                      //      .readdata
		.za_valid       (m_readdatavalid),                 //      .readdatavalid
		.za_waitrequest (m_waitrequest),                   //      .waitrequest
		.zs_addr        (ram_addr),                        //  wire.export
		.zs_ba          (ram_ba),                          //      .export
		.zs_cas_n       (ram_cas_n),                       //      .export
		.zs_cke         (ram_cke),                         //      .export
		.zs_cs_n        (ram_cs_n),                        //      .export
		.zs_dq          (ram_dq),                          //      .export
		.zs_dqm         (ram_dqm),                         //      .export
		.zs_ras_n       (ram_ras_n),                       //      .export
		.zs_we_n        (ram_we_n)                         //      .export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
